--*****************************************************************************
--*  Copyright (c) 2012 by Michael Fischer. All rights reserved.
--*
--*  Redistribution and use in source and binary forms, with or without 
--*  modification, are permitted provided that the following conditions 
--*  are met:
--*  
--*  1. Redistributions of source code must retain the above copyright 
--*     notice, this list of conditions and the following disclaimer.
--*  2. Redistributions in binary form must reproduce the above copyright
--*     notice, this list of conditions and the following disclaimer in the 
--*     documentation and/or other materials provided with the distribution.
--*  3. Neither the name of the author nor the names of its contributors may 
--*     be used to endorse or promote products derived from this software 
--*     without specific prior written permission.
--*
--*  THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS 
--*  "AS IS" AND ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT 
--*  LIMITED TO, THE IMPLIED WARRANTIES OF MERCHANTABILITY AND FITNESS 
--*  FOR A PARTICULAR PURPOSE ARE DISCLAIMED. IN NO EVENT SHALL 
--*  THE COPYRIGHT OWNER OR CONTRIBUTORS BE LIABLE FOR ANY DIRECT, INDIRECT, 
--*  INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES (INCLUDING, 
--*  BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES; LOSS 
--*  OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED 
--*  AND ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, 
--*  OR TORT (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF 
--*  THE USE OF THIS SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF 
--*  SUCH DAMAGE.
--*
--*****************************************************************************
--*  History:
--*
--*  14.07.2011  mifi  First Version
--*****************************************************************************


--*****************************************************************************
--*  DEFINE: Library                                                          *
--*****************************************************************************
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;



--*****************************************************************************
--*  DEFINE: Entity                                                           *
--*****************************************************************************

entity sc_fpga is
   port( 
	      --
         -- Input clock 
         --
         CLOCK_50      : in  std_logic;
			LED_GREEN     : out std_logic_vector(7 downto 0);
         KEY           : in  std_logic_vector(1 downto 0);
         SW            : in  std_logic_vector(3 downto 0);
			RPI           : in  std_logic_vector(3 downto 0);
			SS            : in  std_logic;
			SCLK          : in  std_logic;
			MOSI          : in  std_logic;
			MISO          : in  std_logic
			
       );
end entity sc_fpga;

--*****************************************************************************
--*  DEFINE: Architecture                                                     *
--****************************************************************************

architecture syn of sc_fpga is

   --
   -- Define all components which are included here
   --
	component pll
     port ( 
            inclk0   : in  std_logic  := '0';
            c0       : out std_logic ;
            locked   : out std_logic 
          );
   end component pll;

   --
   -- Define all local signals (like static data) here
   --
   signal el_clk       : std_logic;
   signal pll_locked   : std_logic;
   signal counter_data : std_logic_vector(31 downto 0) := (others => '0');  
	signal saved_sw     : std_logic_vector(3 downto 0) := (others => '0');
   signal SPI_signals  : std_logic_vector(7 downto 0) := (others => '0');
begin

   inst_pll : pll
      port map ( 
                 inclk0 => CLOCK_50,
                 c0     => el_clk,
                 locked => pll_locked
               );

   process(el_clk)
   begin
      if rising_edge(el_clk) then
		  if(SW = saved_sw) then
          counter_data <= std_logic_vector(unsigned(counter_data) + 1);
		  else
			 counter_data <= (others => '0');
		  end if;
		saved_sw <= SW;  
	   end if; 
   end process;
	
  
   SPI_signals(0) <= SS;
	SPI_signals(1) <= MOSI;
	SPI_signals(2) <= MISO;
	SPI_signals(3) <= SCLK;
	
   LED_GREEN <= counter_data(21 downto 14) when saved_sw="0000" else
                SPI_signals                when saved_sw="1111" else
                (others => counter_data(14));
   
end architecture syn;

-- *** EOF ***
